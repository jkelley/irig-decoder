module irig(input         clk_10mhz,
            input         rst,
			input         irigb,
            output        pps,
            output [5:0]  ts_second,
            output [5:0]  ts_minute,
            output [4:0]  ts_hour,
            output [8:0]  ts_day,
            output [6:0]  ts_year,
            output [16:0] ts_sec_day);
    
    wire                  irig_d0;
    wire                  irig_d1;
    wire                  irig_mark;
    wire                  pps_gate;
    wire [3:0]            ts_select;
    wire                  ts_reset;
    wire [3:0]            bit_idx;
    wire [1:0]            digit_idx;
    wire                  bit_value;

    // Decode the IRIG-B width-encoded bits
    // into data 0, data 1, and mark signals
    irig_width_decode id1(.clk(clk_10mhz),
                          .rst(rst),
                          .irigb(irigb),
                          .irig_mark(irig_mark),
                          .irig_d0(irig_d0),
                          .irig_d1(irig_d1));

    // Lock onto and track the IRIG-B "states"
    // separated by mark signals.  Grab the BCD and binary
    // bit values and send them to the timestamp block.
    irig_state is1(.clk(clk_10mhz),
                   .rst(rst),
                   .irig_d0(irig_d0),
                   .irig_d1(irig_d1),
                   .irig_mark(irig_mark),
                   .pps_gate(pps_gate),
                   .ts_select(ts_select),
                   .ts_reset(ts_reset),
                   .bit_idx(bit_idx),
                   .digit_idx(digit_idx),
                   .bit_value(bit_value));

    // From the BCD and binary bit values, generate
    // the timestamps of the previous whole second
    irig_timestamp it1(.clk(clk_10mhz),
                       .rst(rst),
                       .bit_idx(bit_idx),
                       .digit_idx(digit_idx),
                       .bit_value(bit_value),
                       .ts_select(ts_select),
                       .ts_reset(ts_reset),
                       .ts_second(ts_second),
                       .ts_minute(ts_minute),
                       .ts_hour(ts_hour),
                       .ts_day(ts_day),
                       .ts_year(ts_year),
                       .ts_sec_day(ts_sec_day));

    // PPS signal is generated by gating the IRIG signal
    // during the start marker.  Technically this should be a
    // negedge-registered signal, but it is directly
    // generated from the change in the IRIG signal itself
    // so will be set up in time. 
    assign pps = irigb & pps_gate;

endmodule

            
