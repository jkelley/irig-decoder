module irig_timestamp (
	                   input  clk,
                       input  irigb,
	                   input  irig_d0,
	                   input  irig_d1,
	                   input  irig_mark,
	                   output pps,
	                   output reg [16:0] ts_seconds,
	                   input  rst
                       );

    localparam ST_UNLOCKED = 4'd0,
      ST_PRELOCK  = 4'b1,
      ST_START    = 4'd2,
      ST_SECONDS  = 4'd3,
      ST_MINUTES  = 4'd4,
      ST_HOURS    = 4'd5,
      ST_DAYS     = 4'd6,
      ST_DAYS2    = 4'd7,
      ST_YEAR     = 4'd8,
      ST_UNUSED1  = 4'd9,
      ST_UNUSED2  = 4'd10,
      ST_SEC_DAY  = 4'd11,
      ST_SEC_DAY2 = 4'd12;

    // PPS generation
    reg                       pps_en, pps_en_dly;

    // Current and next state machine state
    reg [3:0]                 state, next_state;

    // Count IRIG bits within a state (100/sec)
    reg [3:0]                 irig_cnt;

    // Timestamp generation logic
    reg                       ts_reset;
    reg [16:0]                ts_seconds_mask;

    // PPS signal is generated by gating the IRIG signal
    // during the start marker.  Technically this should be a
    // negedge-registered signal, but it is directly
    // generated from the change in the IRIG signal so should
    // be set up.
    assign pps = irigb & pps_en_dly;

    // Registers
    always @(posedge clk) begin
	    if (rst) begin
		    state <= ST_UNLOCKED;
            pps_en_dly <= 1'b0;
            irig_cnt <= 4'b0;
            ts_seconds <= 17'b0;
        end
	    else begin
		    state <= next_state;
            pps_en_dly <= pps_en;

            // Count the IRIG bits received between every MARK
            if (irig_mark)
              irig_cnt <= 4'b0;
            else 
              irig_cnt <= irig_cnt + (irig_d0 | irig_d1);

            // Reset all the timestamp outputs
            if (ts_reset) begin
                ts_seconds <= 17'b0;
            end
            else begin
                ts_seconds = ts_seconds | ts_seconds_mask;
            end            
        end
    end

    // IRIG decoding state machine
    // FIX ME add timestamp decoding
    always @(*) begin
        next_state = state;
        pps_en = 1'b0;
        ts_reset = 1'b0;
        ts_seconds_mask = 17'b0;
	    case (state)
	      ST_UNLOCKED: begin
		      if (irig_mark)
			    next_state = ST_PRELOCK;
	      end
          ST_PRELOCK: begin
		      if (irig_mark)
			    next_state = ST_SECONDS;
		      else if (irig_d0 || irig_d1)
			    next_state = ST_UNLOCKED;          
          end
	      ST_START: begin
              pps_en = 1'b1;
		      if (irig_mark) begin
                  ts_reset = 1'b1;
				  next_state = ST_SECONDS;
              end
	      end
	      ST_SECONDS: begin
		      if (irig_mark)
			    next_state = ST_MINUTES;
	      end
	      ST_MINUTES: begin
		      if (irig_mark)
			    next_state = ST_HOURS;
	      end		
	      ST_HOURS: begin
		      if (irig_mark)
			    next_state = ST_DAYS;
	      end
	      ST_DAYS: begin
		      if (irig_mark)
			    next_state = ST_DAYS2;
	      end
	      ST_DAYS2: begin
		      if (irig_mark)
			    next_state = ST_YEAR;
	      end
	      ST_YEAR: begin
		      if (irig_mark)
			    next_state = ST_UNUSED1;
	      end
	      ST_UNUSED1: begin
		      if (irig_mark)
			    next_state = ST_UNUSED2;
	      end
	      ST_UNUSED2: begin
		      if (irig_mark)
			    next_state = ST_SEC_DAY;
	      end
	      ST_SEC_DAY: begin
              ts_seconds_mask = irig_d1 << irig_cnt;
		      if (irig_mark)
			    next_state = ST_SEC_DAY2;
	      end
	      ST_SEC_DAY2: begin
              ts_seconds_mask = irig_d1 << (irig_cnt+9);
		      if (irig_mark) begin
			      next_state = ST_START;
                  pps_en = 1'b1;
              end
	      end
	    endcase
    end
    
endmodule
